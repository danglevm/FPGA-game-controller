module ACCELEROMETER
#(
	parameter c_SPI_CLK_FREQ
)
()