module ACCELEROMETER();

endmodule